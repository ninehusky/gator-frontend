module constant (input a, output blah);
    assign blah = 1;
endmodule